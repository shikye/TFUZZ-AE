assign prefix_inst_storage = '{
    64'h11828293_00000297,
    64'h00000093_30529073,
    64'h00000193_00000113,
    64'h00000293_00000213,
    64'h00000393_00000313,
    64'h00000493_00000413,
    64'h00000593_00000513,
    64'h00000693_00000613,
    64'h00000793_00000713,
    64'h00000893_00000813,
    64'h00000993_00000913,
    64'h00000a93_00000a13,
    64'h00000b93_00000b13,
    64'h00000c93_00000c13,
    64'h00000d93_00000d13,
    64'h00000e93_00000e13,
    64'h00000f93_00000f13,
    64'h30052073_00006537,
    64'hf2000053_00305073,
    64'hf2000153_f20000d3,
    64'hf2000253_f20001d3,
    64'hf2000353_f20002d3,
    64'hf2000453_f20003d3,
    64'hf2000553_f20004d3,
    64'hf2000653_f20005d3,
    64'hf2000753_f20006d3,
    64'hf2000853_f20007d3,
    64'hf2000953_f20008d3,
    64'hf2000a53_f20009d3,
    64'hf2000b53_f2000ad3,
    64'hf2000c53_f2000bd3,
    64'hf2000d53_f2000cd3,
    64'hf2000e53_f2000dd3,
    64'hf2000f53_f2000ed3,
    64'h0440006f_f2000fd3,
    64'h00200313_342022f3,
    64'h00000033_00530863,
    64'h00000033_00000033,
    64'h00d2d293_300022f3,
    64'h00028863_0032f293,
    64'h00000033_00000033,
    64'h00006537_00000033,
    64'h30200073_30052073
};

// Total bytes: 344
